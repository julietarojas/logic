//: version "2.0-b10"
//: property encoding = "iso8859-1"
//: property locale = "en"
//: property prefix = "_GG"
//: property title = "subtractor.v"
//: property timingViolationMode = 2
//: property initTime = "0 ns"

`timescale 1ns/1ns

//: /netlistBegin main
module main;    //: root_module
reg [7:0] B;    //: /sn:0 {0}(#:366,163)(366,262)(421,262)(421,277){1}
reg [7:0] A;    //: /sn:0 {0}(#:507,163)(507,262)(453,262)(453,277){1}
reg w1;    //: /sn:0 {0}(405,339)(405,332)(334,332){1}
supply0 w5;    //: /sn:0 {0}(461,291)(470,291){1}
//: {2}(474,291)(491,291)(491,317){3}
//: {4}(472,293)(472,353)(445,353){5}
wire [7:0] w6;    //: /sn:0 {0}(#:656,311)(656,383){1}
//: {2}(#:654,385)(550,385)(550,245){3}
//: {4}(656,387)(656,444)(421,444)(421,401){5}
//: {6}(421,400)(#:421,368){7}
wire w4;    //: /sn:0 {0}(413,291)(398,291){1}
wire w3;    //: /sn:0 {0}(425,401)(613,401)(613,292)(604,292){1}
wire w8;    //: /sn:0 {0}(397,353)(382,353){1}
wire [7:0] w2;    //: /sn:0 {0}(#:437,306)(437,339){1}
//: enddecls

  //: joint g4 (w5) @(472, 291) /w:[ 2 -1 1 4 ]
  _GGADD8 #(68, 70, 62, 64) g8 (.A(w1), .B(w2), .S(w6), .CI(w5), .CO(w8));   //: @(421,355) /sn:0 /w:[ 0 1 7 5 0 ]
  //: LED g3 (w3) @(597,292) /sn:0 /R:1 /w:[ 1 ] /type:0
  //: GROUND g2 (w5) @(491,323) /sn:0 /w:[ 3 ]
  //: LED g1 (w6) @(656,304) /sn:0 /w:[ 0 ] /type:3
  //: LED g11 (w6) @(550,238) /sn:0 /w:[ 3 ] /type:2
  //: SWITCH g10 (w1) @(317,332) /sn:0 /w:[ 1 ] /st:0 /dn:1
  //: DIP g6 (A) @(507,153) /sn:0 /w:[ 0 ] /st:0 /dn:1
  assign w3 = w6[7]; //: TAP g9 @(419,401) /sn:0 /R:2 /w:[ 0 5 6 ] /ss:1
  //: comment g7 @(334,333) /sn:0
  //: /line:"<b>signo<b>"
  //: /end
  //: DIP g5 (B) @(366,153) /sn:0 /w:[ 0 ] /st:0 /dn:1
  _GGADD8 #(70, 72, 62, 64) g0 (.A(~B), .B(A), .S(w2), .CI(w5), .CO(w4));   //: @(437,293) /sn:0 /w:[ 1 1 0 0 0 ]
  //: joint g12 (w6) @(656, 385) /w:[ -1 1 2 4 ]

endmodule
//: /netlistEnd
