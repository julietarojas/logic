//: version "2.0-b10"
//: property encoding = "iso8859-1"
//: property locale = "en"
//: property prefix = "_GG"
//: property timingViolationMode = 2
//: property initTime = "0 ns"

`timescale 1ns/1ns

//: /netlistBegin main
module main;    //: root_module
reg w0;    //: /sn:0 {0}(212,77)(183,77)(183,77)(156,77){1}
reg w1;    //: /sn:0 {0}(212,271)(181,271)(181,271)(149,271){1}
wire w6;    //: /sn:0 {0}(233,274)(263,274)(263,245)(269,245){1}
wire w7;    //: /sn:0 {0}(290,243)(319,243){1}
//: {2}(323,243)(351,243)(351,216){3}
//: {4}(321,241)(321,109)(266,109)(266,94)(276,94){5}
wire w4;    //: /sn:0 {0}(233,80)(259,80)(259,89)(276,89){1}
wire w3;    //: /sn:0 {0}(145,307)(197,307)(197,278){1}
//: {2}(199,276)(212,276){3}
//: {4}(197,274)(197,82)(212,82){5}
wire w8;    //: /sn:0 {0}(339,63)(339,92)(330,92){1}
//: {2}(326,92)(297,92){3}
//: {4}(328,94)(328,225)(259,225)(259,240)(269,240){5}
//: enddecls

  //: joint g8 (w7) @(321, 243) /w:[ 2 4 1 -1 ]
  _GGNAND2 #(4) g4 (.I0(w4), .I1(w7), .Z(w8));   //: @(287,92) /sn:0 /w:[ 1 5 3 ]
  _GGNAND2 #(4) g3 (.I0(w1), .I1(w3), .Z(w6));   //: @(223,274) /sn:0 /w:[ 0 3 0 ]
  _GGNAND2 #(4) g2 (.I0(w0), .I1(w3), .Z(w4));   //: @(223,80) /sn:0 /w:[ 0 5 0 ]
  //: SWITCH g1 (w1) @(132,271) /sn:0 /w:[ 1 ] /st:0 /dn:1
  //: joint g11 (w3) @(197, 276) /w:[ 2 4 -1 1 ]
  _GGCLOCK_P100_0_50 g10 (.Z(w3));   //: @(132,307) /sn:0 /w:[ 0 ] /omega:100 /phi:0 /duty:50
  //: LED g6 (w8) @(339,56) /sn:0 /w:[ 0 ] /type:0
  //: joint g9 (w8) @(328, 92) /w:[ 1 -1 2 4 ]
  //: LED g7 (w7) @(351,209) /sn:0 /w:[ 3 ] /type:0
  _GGNAND2 #(4) g5 (.I0(w8), .I1(w6), .Z(w7));   //: @(280,243) /sn:0 /w:[ 5 1 0 ]
  //: SWITCH g0 (w0) @(139,77) /sn:0 /w:[ 1 ] /st:0 /dn:1

endmodule
//: /netlistEnd
