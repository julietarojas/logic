//: property prefix = "_GG"
//: property title = "BitAdder.v"
//: property timingViolationMode = 2
//: property initTime = "0 ns"

`timescale 1ns/1ns

//: /netlistBegin main
module main;    //: root_module
reg [3:0] B;    //: /sn:0 {0}(#:840,-120)(840,-105){1}
reg [3:0] A;    //: /sn:0 {0}(#:975,-82)(975,-62){1}
//: {2}(975,-61)(975,-44){3}
//: {4}(975,-43)(975,-26){5}
//: {6}(975,-25)(975,5){7}
//: {8}(975,6)(975,18){9}
reg a1;    //: /sn:0 {0}(99,138)(99,161)(170,161){1}
reg b1;    //: /sn:0 {0}(72,177)(170,177){1}
reg a0;    //: /sn:0 {0}(131,51)(131,88)(169,88){1}
reg b0;    //: /sn:0 {0}(61,70)(61,104)(169,104){1}
supply0 w9;    //: /sn:0 {0}(1196,69)(1196,66)(1163,66)(1163,81){1}
wire w6;    //: /sn:0 {0}(288,177)(424,177)(424,53){1}
wire w7;    //: /sn:0 {0}(288,161)(393,161)(393,54){1}
wire w16;    //: /sn:0 {0}(970,-43)(740,-43)(740,64){1}
wire w14;    //: /sn:0 {0}(708,-81)(708,47)(724,47)(724,64){1}
wire w19;    //: /sn:0 {0}(1229,198)(1229,211)(1064,211)(1064,58)(1048,58)(1048,65){1}
wire w4;    //: /sn:0 {0}(970,-61)(899,-61)(899,65){1}
wire w0;    //: /sn:0 {0}(834,186)(834,199)(854,199)(854,55)(867,55)(867,65){1}
wire w3;    //: /sn:0 {0}(287,88)(327,88)(327,56){1}
wire w21;    //: /sn:0 {0}(979,-25)(1080,-25)(1080,65){1}
wire w23;    //: /sn:0 {0}(832,185)(1080,185)(1080,179){1}
wire w20;    //: /sn:0 {0}(728,-81)(728,50)(1064,50)(1064,65){1}
wire w1;    //: /sn:0 {0}(718,-81)(718,51)(883,51)(883,65){1}
wire w25;    //: /sn:0 {0}(738,-81)(738,54)(1212,54)(1212,69){1}
wire w18;    //: /sn:0 {0}(740,178)(740,208)(741,208)(741,223){1}
wire w8;    //: /sn:0 {0}(708,64)(708,54)(723,54)(723,83)(884,83)(884,189)(899,189)(899,179){1}
wire w22;    //: /sn:0 {0}(1064,179)(1064,199)(1064,199)(1064,222){1}
wire w17;    //: /sn:0 {0}(724,178)(724,203)(724,203)(724,222){1}
wire [1:0] w12;    //: /sn:0 {0}(#:723,-87)(723,-106)(838,-106){1}
wire w2;    //: /sn:0 {0}(287,104)(356,104)(356,55){1}
wire w27;    //: /sn:0 {0}(1212,183)(1212,197)(1212,197)(1212,222){1}
wire w5;    //: /sn:0 {0}(883,179)(883,203)(883,203)(883,222){1}
wire w29;    //: /sn:0 {0}(1228,198)(1228,183){1}
wire w26;    //: /sn:0 {0}(979,6)(1228,6)(1228,69){1}
//: enddecls

  //: LED g8 (w2) @(356,48) /sn:0 /w:[ 1 ] /type:0
  //: SWITCH g4 (a1) @(99,125) /sn:0 /R:3 /w:[ 0 ] /st:0 /dn:1
  sumador g13 (.a(w21), .b(w20), .cin(w19), .cout(w23), .s(w22));   //: @(1032, 66) /sz:(64, 112) /R:3 /sn:0 /p:[ Ti0>1 Ti1>1 Ti2>1 Bo0<1 Bo1<0 ]
  //: SWITCH g3 (b0) @(61,57) /sn:0 /R:3 /w:[ 0 ] /st:0 /dn:1
  //: SWITCH g2 (a0) @(131,38) /sn:0 /R:3 /w:[ 0 ] /st:0 /dn:1
  semisumador g1 (.a0(a1), .b0(b1), .c(w7), .s0(w6));   //: @(171, 145) /sz:(116, 48) /sn:0 /p:[ Li0>1 Li1>1 Ro0<0 Ro1<0 ]
  //: DIP g11 (B) @(840,-130) /sn:0 /w:[ 0 ] /st:0 /dn:1
  //: DIP g16 (A) @(975,-92) /sn:0 /w:[ 0 ] /st:0 /dn:1
  sumador g10 (.a(w4), .b(w1), .cin(w0), .cout(w8), .s(w5));   //: @(851, 66) /sz:(64, 112) /R:3 /sn:0 /p:[ Ti0>1 Ti1>1 Ti2>1 Bo0<1 Bo1<0 ]
  //: LED g27 (w18) @(741,230) /sn:0 /R:2 /w:[ 1 ] /type:0
  assign w4 = A[2]; //: TAP g19 @(973,-61) /sn:0 /R:2 /w:[ 0 2 1 ] /ss:0
  //: LED g6 (w3) @(327,49) /sn:0 /w:[ 1 ] /type:0
  //: LED g9 (w6) @(424,46) /sn:0 /w:[ 1 ] /type:0
  //: LED g7 (w7) @(393,47) /sn:0 /w:[ 1 ] /type:0
  assign w16 = A[3]; //: TAP g20 @(973,-43) /sn:0 /R:2 /w:[ 0 4 3 ] /ss:0
  //: LED g15 (w27) @(1212,229) /sn:0 /R:2 /w:[ 1 ] /type:0
  //: LED g25 (w5) @(883,229) /sn:0 /R:2 /w:[ 1 ] /type:0
  assign w26 = A[0]; //: TAP g17 @(973,6) /sn:0 /R:2 /w:[ 0 8 7 ] /ss:1
  sumador g14 (.a(w26), .b(w25), .cin(w9), .cout(w29), .s(w27));   //: @(1180, 70) /sz:(64, 112) /R:3 /sn:0 /p:[ Ti0>1 Ti1>1 Ti2>0 Bo0<1 Bo1<0 ]
  //: SWITCH g5 (b1) @(55,177) /sn:0 /w:[ 0 ] /st:0 /dn:1
  //: LED g24 (w17) @(724,229) /sn:0 /R:2 /w:[ 1 ] /type:0
  //: GROUND g21 (w9) @(1163,87) /sn:0 /w:[ 1 ]
  //: LED g26 (w22) @(1064,229) /sn:0 /R:2 /w:[ 1 ] /type:0
  tran g22[1:0] ({w25, w20, w1, w14}, w12);   //: @(723,-86) /sn:0 /R:1 /dr:0 /tp:0 /drp:-1 /w:[ 0 0 0 0 0 ]
  semisumador g0 (.a0(a0), .b0(b0), .c(w3), .s0(w2));   //: @(170, 72) /sz:(116, 48) /sn:0 /p:[ Li0>1 Li1>1 Ro0<0 Ro1<0 ]
  assign w21 = A[1]; //: TAP g18 @(973,-25) /sn:0 /R:2 /w:[ 0 6 5 ] /ss:1
  sumador g12 (.a(w16), .b(w14), .cin(w8), .cout(w18), .s(w17));   //: @(692, 65) /sz:(64, 112) /R:3 /sn:0 /p:[ Ti0>1 Ti1>1 Ti2>0 Bo0<0 Bo1<0 ]

endmodule
//: /netlistEnd

//: /netlistBegin sumador
module sumador(s, b, a, cout, cin);
//: interface  /sz:(112, 64) /bd:[ Li0>cin(48/64) Li1>b(32/64) Li2>a(16/64) Ro0<s(32/64) Ro1<cout(16/64) ] /pd: 0 /pi: 0 /pe: 1 /pp: 1
input b;    //: /sn:0 {0}(158,203)(185,203){1}
//: {2}(189,203)(363,203)(363,118)(371,118){3}
//: {4}(187,201)(187,183)(239,183){5}
//: {6}(187,205)(187,226)(240,226){7}
input cin;    //: /sn:0 {0}(169,108)(197,108){1}
//: {2}(201,108)(371,108){3}
//: {4}(199,110)(199,130){5}
//: {6}(201,132)(238,132){7}
//: {8}(199,134)(199,178)(239,178){9}
output s;    //: /sn:0 {0}(392,113)(445,113){1}
input a;    //: /sn:0 {0}(160,149)(205,149){1}
//: {2}(209,149)(319,149)(319,113)(371,113){3}
//: {4}(207,151)(207,221)(240,221){5}
output cout;    //: /sn:0 {0}(315,181)(398,181){1}
wire w3;    //: /sn:0 {0}(294,186)(276,186)(276,224)(261,224){1}
wire w0;    //: /sn:0 {0}(294,176)(273,176)(273,135)(259,135){1}
wire w1;    //: /sn:0 {0}(294,181)(260,181){1}
wire w10;    //: /sn:0 {0}(207,168)(218,168){1}
//: {2}(220,166)(220,137)(238,137){3}
//: {4}(220,170)(220,172){5}
//: enddecls

  _GGAND2 #(6) g8 (.I0(cin), .I1(b), .Z(w1));   //: @(250,181) /sn:0 /w:[ 9 5 1 ]
  //: OUT g4 (s) @(442,113) /sn:0 /w:[ 1 ]
  //: joint g13 (b) @(187, 203) /w:[ 2 4 1 6 ]
  _GGXOR3 #(11) g3 (.I0(cin), .I1(a), .I2(b), .Z(s));   //: @(382,113) /sn:0 /w:[ 3 3 3 0 ]
  //: IN g2 (b) @(156,203) /sn:0 /w:[ 0 ]
  //: IN g1 (a) @(158,149) /sn:0 /w:[ 0 ]
  //: joint g11 (cin) @(199, 132) /w:[ 6 5 -1 8 ]
  //: joint g10 (cin) @(199, 108) /w:[ 2 -1 1 4 ]
  //: OUT g6 (cout) @(395,181) /sn:0 /w:[ 1 ]
  _GGAND2 #(6) g9 (.I0(cin), .I1(w10), .Z(w0));   //: @(249,135) /sn:0 /w:[ 7 3 1 ]
  _GGAND2 #(6) g7 (.I0(a), .I1(b), .Z(w3));   //: @(251,224) /sn:0 /w:[ 5 7 1 ]
  //: joint g14 (w10) @(220, 168) /w:[ -1 2 1 4 ]
  _GGOR3 #(8) g5 (.I0(w0), .I1(w1), .I2(w3), .Z(cout));   //: @(305,181) /sn:0 /w:[ 0 0 0 0 ]
  //: IN g0 (cin) @(167,108) /sn:0 /w:[ 0 ]
  //: joint g12 (a) @(207, 149) /w:[ 2 -1 1 4 ]

endmodule
//: /netlistEnd

//: /netlistBegin semisumador
module semisumador(c, s0, b0, a0);
//: interface  /sz:(116, 48) /bd:[ Li0>b0(32/48) Li1>a0(16/48) Ro0<s0(32/48) Ro1<c(16/48) ] /pd: 0 /pi: 0 /pe: 1 /pp: 1
output s0;    //: /sn:0 {0}(236,44)(160,44){1}
input a0;    //: /sn:0 {0}(-2,43)(36,43){1}
//: {2}(40,43)(43,43)(43,98)(56,98){3}
//: {4}(38,41)(38,26)(63,26){5}
input b0;    //: /sn:0 {0}(2,112)(16,112){1}
//: {2}(20,112)(43,112)(43,103)(56,103){3}
//: {4}(18,110)(18,61){5}
//: {6}(20,59)(62,59){7}
//: {8}(18,57)(18,31)(63,31){9}
output c;    //: /sn:0 {0}(176,101)(77,101){1}
wire w7;    //: /sn:0 {0}(5,43)(5,54)(62,54){1}
wire w0;    //: /sn:0 {0}(84,29)(124,29)(124,41)(139,41){1}
wire w1;    //: /sn:0 {0}(83,57)(124,57)(124,46)(139,46){1}
//: enddecls

  //: joint g8 (b0) @(18, 112) /w:[ 2 4 1 -1 ]
  _GGAND2 #(6) g4 (.I0(a0), .I1(b0), .Z(c));   //: @(67,101) /sn:0 /w:[ 3 3 1 ]
  //: OUT g3 (c) @(173,101) /sn:0 /w:[ 0 ]
  //: OUT g2 (s0) @(233,44) /sn:0 /w:[ 0 ]
  //: IN g1 (b0) @(0,112) /sn:0 /w:[ 0 ]
  //: joint g10 (a0) @(38, 43) /w:[ 2 4 1 -1 ]
  _GGAND2 #(6) g6 (.I0(a0), .I1(!b0), .Z(w0));   //: @(74,29) /sn:0 /w:[ 5 9 0 ]
  //: joint g9 (b0) @(18, 59) /w:[ 6 8 -1 5 ]
  _GGAND2 #(6) g7 (.I0(!w7), .I1(b0), .Z(w1));   //: @(73,57) /sn:0 /w:[ 1 7 0 ]
  _GGOR2 #(6) g5 (.I0(w0), .I1(w1), .Z(s0));   //: @(150,44) /sn:0 /w:[ 1 1 1 ]
  //: IN g0 (a0) @(-4,43) /sn:0 /w:[ 0 ]

endmodule
//: /netlistEnd
